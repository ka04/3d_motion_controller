`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   23:22:07 04/08/2014
// Design Name:   CF
// Module Name:   C:/Users/YangTianyu/Desktop/EC551/CompFilter/TB_CF.v
// Project Name:  CompFilter
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: CF
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module TB_CF;

	// Inputs
	reg [15:0] gyroData;
	reg [15:0] y_accel_data;
	reg [15:0] z_accel_data;
	reg clk;
	reg RST;

	// Outputs
	wire [15:0] x_temp;
	wire [31:0] x_final;

	// Instantiate the Unit Under Test (UUT)
	CF uut (
		.gyroData(gyroData), 
		.y_accel_data(y_accel_data), 
		.z_accel_data(z_accel_data), 
		.clk(clk), 
		.RST(RST),
		.x_temp(x_temp), 
		.x_final(x_final)
	);

	initial begin
		clk = 0;RST=0;
		// Initialize Inputs
		
		#50 RST=1; gyroData = 16'h0080;y_accel_data = 16'h1000;z_accel_data = 16'h1000;
		#50 gyroData = 16'h0100;y_accel_data = 16'h1000;z_accel_data = 16'h1000;
		#50 gyroData = 16'h0200;y_accel_data = 16'h1000;z_accel_data = 16'h2000;
		#50 gyroData = 16'h0400;y_accel_data = 16'h1000;z_accel_data = 16'h3000;
		#50 gyroData = 16'h0800;y_accel_data = 16'h1000;z_accel_data = 16'h4000;


		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here
	end
      
		always begin
		#10 clk = ~clk;
		end
		
		
		
endmodule

